library verilog;
use verilog.vl_types.all;
entity Timer_tb is
end Timer_tb;
